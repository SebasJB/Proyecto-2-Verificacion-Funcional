class c_1882_4;
    bit[31:0] seq_id = 32'he;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1882_4;
    c_1882_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxx0110xzzx0z0xxz1z101x0xz0zz11xxzzzzxxzxxzzzzzzxxzxzzxxzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
