class c_975_4;
    bit[31:0] seq_id = 32'h2;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_975_4;
    c_975_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10x0x1x1zx0xzxxz1x1zz1zz0x10z1xzzzzzzxzxxxxxzxxxzzzxzzzzxxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
