class c_1342_4;
    bit[31:0] seq_id = 32'h8;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1342_4;
    c_1342_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxxxz00z1zzx10z1z1z1z1x101xx10zxxxxxxzxzxzxzzxxxzxzzzzzzzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
