class c_81_4;
    bit[31:0] seq_id = 32'h9;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_81_4;
    c_81_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x00x111x1xxz1101z1x0z0z00z0x101zxzzzzzzzxzxzzzxxxzxzzxzzxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
