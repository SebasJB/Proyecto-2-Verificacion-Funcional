class c_1402_4;
    bit[31:0] seq_id = 32'h4;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1402_4;
    c_1402_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10101x11z1011x11x1z11z1z00x1110xzxzxxzxzxzzzxzxzxxzxxzxxzxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
