class c_1363_4;
    bit[31:0] seq_id = 32'h2;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1363_4;
    c_1363_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10x0z00zxzz1x0x1x100z1zz0z0zxzx1xzzxzxzxzzxxxzxxzzxxxxzzzzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
