class c_968_4;
    bit[31:0] seq_id = 32'h9;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_968_4;
    c_968_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zx11z1z1xz0xzzx1x1z000x11xzzx1zzxxzxxzzxzzxzxxxxxxxzxxxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
