class c_1860_4;
    bit[31:0] seq_id = 32'h7;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1860_4;
    c_1860_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xx00z00zxxx1xzxz0z0110z01z1z10zzzzzzxxzzxxzzxzxxzxxzzxzzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
