class c_457_4;
    bit[31:0] seq_id = 32'hf;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_457_4;
    c_457_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x011xxx1xx1zxzzxzz00zzx01010xxxzxxzxxzzxzzxxzzzxxxzxzzxxxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
