class c_1889_4;
    bit[31:0] seq_id = 32'ha;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1889_4;
    c_1889_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx01xzxzx1zzx0zx00010z0x1x10xz0zxzxzxzxzzxzxxzzzxxzxzxxzxzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
