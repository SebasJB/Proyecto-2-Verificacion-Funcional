class c_28_4;
    bit[31:0] seq_id = 32'hc;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_28_4;
    c_28_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111x1zzx00x1z1x0x001xxx001zxzxzxzxxzxxzzxxzzzzzzzxxzzzzzxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
