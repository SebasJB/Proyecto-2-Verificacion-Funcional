class c_64_4;
    bit[31:0] seq_id = 32'h0;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_64_4;
    c_64_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxxzx1z000z0zz1xzz1z0x00x1xz00xxzxzzzxxzzzzzzzxxxzxzxxxxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
