class c_99_4;
    bit[31:0] seq_id = 32'ha;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_99_4;
    c_99_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11z0x1x0x0xz1x1xz01xx1xx1zx0100xzxxzzzxxzzxxzzxzzxzxzzzxzxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
