class c_1415_4;
    bit[31:0] seq_id = 32'he;
    bit[7:0] pkt_id = 8'h0;
    integer t = 3;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1415_4;
    c_1415_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxzxx11z0x101z0z10z0z01xx1x1xz1zxzzzxxzzzzxxzzzzzxxxxzxxxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
