class c_119_4;
    bit[31:0] seq_id = 32'h3;
    bit[7:0] pkt_id = 8'h0;
    integer t = 3;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_119_4;
    c_119_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z01x1x0x01x1zxz10xx1zzxx0z1x01zxxzxzxzzxxxzxzxzzxzxzxzzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
