class c_1857_4;
    bit[31:0] seq_id = 32'ha;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1857_4;
    c_1857_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z1x01xx11x0z1zx1x110001x11xxx0zxzzxxxzxzxzxzzxxzxxzzxxzxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
