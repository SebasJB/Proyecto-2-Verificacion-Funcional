class c_59_4;
    bit[31:0] seq_id = 32'hd;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_59_4;
    c_59_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xzx00xz11z10zzzxxx00zxzx1x010zxxzzzzxxzxzxxzzzzxzxxxzzzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
