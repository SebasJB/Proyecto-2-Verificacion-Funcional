class c_462_4;
    bit[31:0] seq_id = 32'ha;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_462_4;
    c_462_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10z111z0xxx0z0x1zx01zzzz0110z1zxxxzzzxzzzxxzxxxzxxxxxzzzxxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
