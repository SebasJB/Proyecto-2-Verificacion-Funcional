class c_1872_4;
    bit[31:0] seq_id = 32'h4;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1872_4;
    c_1872_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1xx01z10zzz1x1xz1xx00z0zxxzz0xxzzxxxzxxzxxzzzxxxzzxxxzxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
