class c_1357_4;
    bit[31:0] seq_id = 32'h8;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1357_4;
    c_1357_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0x1zzx0001zzzxz1z01xzx0z1100x1zxxxxxzxxxxxxzxzxzxzxzxxxzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
