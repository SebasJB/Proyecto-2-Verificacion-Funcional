class c_1903_4;
    bit[31:0] seq_id = 32'h3;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1903_4;
    c_1903_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0xz001x0x0xx0x00xzxz11zx000zzxxxzzxzxxzzxxxzxxzxzxxxzzzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
