class c_1899_4;
    bit[31:0] seq_id = 32'h0;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1899_4;
    c_1899_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zzxz11zz111x0010z101x1zx1x0x10xzzxzxxzzxxxzxxxzzxxzxzzxzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
