class c_1029_4;
    bit[31:0] seq_id = 32'hc;
    bit[7:0] pkt_id = 8'h0;
    integer t = 3;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1029_4;
    c_1029_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11z01xzx0x11z0zzxx0x00zxxzz1111xxzxzzxxxxzxxzzzzxzzxzxxzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
