class c_1320_4;
    bit[31:0] seq_id = 32'hd;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1320_4;
    c_1320_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1z0x0z00x10z11zx01zzx0101z1xxxxzzxzxxxxzxzxzxzxxzxzxxxxzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
