class c_448_4;
    bit[31:0] seq_id = 32'h7;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_448_4;
    c_448_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z0011xx0zz111x1x0z010x0z100z00zzzzxxzzxxxzzzxxxxxxzzxxxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
