class c_953_4;
    bit[31:0] seq_id = 32'h7;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_953_4;
    c_953_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx0x111001zzx10xx0000x01x1zx11xzxxzxxzzxxxxzxxzzxxxzzzzxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
