class c_26_4;
    bit[31:0] seq_id = 32'he;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_26_4;
    c_26_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1zx1xxxz0z1x1xz110z011z010x111zxxzxzzzzzxzzxxzxxxzxxzzzxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
