class c_58_4;
    bit[31:0] seq_id = 32'he;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_58_4;
    c_58_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxx0xx01zzxz000x0110zz1zz1z01xxzzxzxxzzzzzzzxzzzzzzxzzxzzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
