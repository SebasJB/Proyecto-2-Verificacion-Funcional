class c_1035_4;
    bit[31:0] seq_id = 32'h6;
    bit[7:0] pkt_id = 8'h0;
    integer t = 3;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1035_4;
    c_1035_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx1zxz0zx1x0z0x00zx0x01z1101zx0zzzxxzxzzzxxzxxxxxzzxzzxzzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
