class c_1019_4;
    bit[31:0] seq_id = 32'h9;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1019_4;
    c_1019_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1011z1x1x1x1zzxz0xzx00zxz0zz1z1zxxzzzzxzzxxzzzxzxzxxzxzxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
