class c_491_4;
    bit[31:0] seq_id = 32'hd;
    bit[7:0] pkt_id = 8'h0;
    integer t = 3;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_491_4;
    c_491_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0111zz01x1x1000zxxz0x1zx1x11x0zzzxzxzzxzzzzzzzzzxzzxzzxxxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
