class c_940_4;
    bit[31:0] seq_id = 32'h5;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_940_4;
    c_940_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zx1z0xzzxxxxz010000zz0x0xz110zxxzxxzxzxzxzzzzzxzzxzzzxxxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
