class c_1025_4;
    bit[31:0] seq_id = 32'hf;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1025_4;
    c_1025_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11xzxx1zxx0x00zz1zzx01xzx0xz1z1xzxxzxxzxzzxzxzzzxzzzxxzxzxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
