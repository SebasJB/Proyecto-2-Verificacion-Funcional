class c_67_4;
    bit[31:0] seq_id = 32'ha;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_67_4;
    c_67_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz00100xzz0xz111x1zxzz0xzz1x11x1zzzzzxxzxzzzxzxxzxzzxxzxxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
