class c_1894_4;
    bit[31:0] seq_id = 32'h5;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1894_4;
    c_1894_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxz0000100zz000z1xx10x000111zz1zxxxzxzzzzxzxxxxxxzzzxxxzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
