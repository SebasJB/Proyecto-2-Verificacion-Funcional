class c_1074_4;
    integer test_mode = 0; // ( test_mode = $unit::scenario_t::GENERAL ) 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:95)
    {
       (test_mode == 1 /* $unit::scenario_t::SATURATION */);
    }
endclass

program p_1074_4;
    c_1074_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1x11z000xxxzxx011zz01zz11x11z0zzxzzzxxzxxxxzzxzzxxxxxzzzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
