class c_464_2;
    bit[4:0] src_id = 5'h0;
    bit[31:0] targets_2_ = 32'h0;
    rand bit[31:0] dest_addr; // rand_mode = ON 

    constraint c_dest_addr_this    // (constraint_mode = ON) (TypesandTransactions.sv:116)
    {
       (dest_addr != src_id);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (dest_addr == targets_2_);
    }
endclass

program p_464_2;
    c_464_2 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10111z0xz1z11z010z10x0z0z0x0111zzzzzzxzzxzzxzxxxxzxzzzzzzxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
