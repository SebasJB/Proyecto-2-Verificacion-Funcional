class c_1914_4;
    bit[31:0] seq_id = 32'he;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1914_4;
    c_1914_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1010zxxzx1011xxzzx0x000010x1x1z1zxzzxzzxzxxzxzxxxxzzxzxxzxxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
