class c_418_4;
    bit[31:0] seq_id = 32'h9;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_418_4;
    c_418_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z0x1xz1z01x1z11xzx1xx1x11zzzz0xxxzxzzxxzxxxzzxxzxxxzxzxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
