class c_446_4;
    bit[31:0] seq_id = 32'h5;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_446_4;
    c_446_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x1xx00xxzx0110z0z1x100111z101z1zzxzzzzxzzxzzzzxzzxzxzzxzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
