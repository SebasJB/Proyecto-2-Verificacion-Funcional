class c_46_4;
    bit[31:0] seq_id = 32'h7;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_46_4;
    c_46_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz101z0z0zz0xx1x01x1x1xz0zz1xz0xxzxzzxzxxxzxzxzxzzzxxzzxzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
