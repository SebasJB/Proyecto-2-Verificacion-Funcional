class c_40_4;
    bit[31:0] seq_id = 32'hf;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_40_4;
    c_40_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0110z1x00x1z101z0zxz01z01xx0x0x1zxxxzxzxxxxzzxzxxxxzzzxzzxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
