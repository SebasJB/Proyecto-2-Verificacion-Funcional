class c_92_4;
    bit[31:0] seq_id = 32'hc;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_92_4;
    c_92_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110xx1zxzzzx1z0zzz10110z0zx11010zxxzzzzzxzxzxxzxxzzzzzzzzxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
