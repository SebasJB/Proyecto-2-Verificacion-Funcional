class c_74_4;
    bit[31:0] seq_id = 32'h3;
    bit[7:0] pkt_id = 8'h0;
    integer t = 1;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_74_4;
    c_74_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x0xxx01z1x11xz0z0zx11x0z00x1xxzzxzzxzxzxxzxxxzzzzxxzzzzxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
