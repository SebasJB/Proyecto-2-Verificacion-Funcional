class c_1858_4;
    bit[31:0] seq_id = 32'h9;
    bit[7:0] pkt_id = 8'h0;
    integer t = 0;
    integer mm = 0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1858_4;
    c_1858_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01xxz0xx0z1xx0z01101z1zzxxzz1x1zzzzxxxzzxxzzxzxxxxxzzxxzxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
