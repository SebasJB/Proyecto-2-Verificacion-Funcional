class c_109_4;
    bit[31:0] seq_id = 32'h6;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_109_4;
    c_109_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx11zx0x01zx1zzzzz0x00x0x1xxx000zxxzzzzxxzzzzzzzxzxzzxxzxzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
