class c_1442_4;
    bit[31:0] seq_id = 32'hc;
    bit[7:0] pkt_id = 8'h0;
    integer t = 3;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1442_4;
    c_1442_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzzz1x00xz1xx1zz1z0zz111zz110xxzxxxxxzxxxxzzxzxxzxzzxxxzxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
