class c_1044_4;
    bit[31:0] seq_id = 32'h2;
    bit[7:0] pkt_id = 8'h0;
    integer t = 3;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1044_4;
    c_1044_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0x0zz101xx1zz10zx001zxx100zz0xxzzxxzzzzzzzxxzzzxzzzxxzzzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
