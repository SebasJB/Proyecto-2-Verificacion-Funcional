class c_1401_4;
    bit[31:0] seq_id = 32'h3;
    bit[7:0] pkt_id = 8'h0;
    integer t = 2;
    integer mm = 1;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (Secuencer.sv:60)
    {
       (pkt_id == (((16 * seq_id) + (t * 2)) + mm));
    }
endclass

program p_1401_4;
    c_1401_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01010zz0x0zzxzzz00zx01xx101zzzzxzzzzxxxzzxzzzxzxzxzxzxxxxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
